ENTITY conte_ate_5 IS
PORT (IN_CLK, RESET: IN BIT;
SAIDA: OUT INTEGER RANGE 0 TO 5;
C_OUT: OUT BIT);
END conte_ate_5;

ARCHITECTURE MASTER OF conte_ate_5 IS
SIGNAL AUX_01: BIT;
SIGNAL AUX_02: INTEGER RANGE 0 TO 5;
BEGIN
PROCESS(IN_CLK)
BEGIN
IF RESET='1' THEN
AUX_02<=0;
AUX_01<='0';
ELSIF (IN_CLK'EVENT)AND(IN_CLK='1')THEN
	IF AUX_02=5 THEN
	AUX_02<=0;
   AUX_01<='1';
	ELSE
	AUX_01<='0';
	AUX_02<=AUX_02+1;
	END IF;
END IF;
END PROCESS;
SAIDA<= AUX_02;
C_OUT<=AUX_01;
END MASTER;			  