ENTITY PRINCIPAL IS
PORT(CLK: IN BIT;
SAI_C1, SAI_C2, SAI_C3: OUT BIT;
ENT_S1, ENT_S2: IN BIT;
DISPLAY_0: OUT BIT_VECTOR ( 6 DOWNTO 0));
END PRINCIPAL;

ARCHITECTURE ONE OF PRINCIPAL IS 
SIGNAL AUX_CLK_TO_FSM: BIT;
SIGNAL AUX_FMS_TO_DEC: INTEGER RANGE 0 TO 7;

COMPONENT DIV_CLK IS
PORT(IN_CLK: IN BIT;
OUT_CLK: OUT BIT);
END COMPONENT;

COMPONENT FMS_ESTPROJ IS
PORT(IN_CLK,S1,S2: IN BIT;
C1, C2, C3: OUT BIT;
DISPLAY_7_SEG: OUT INTEGER RANGE 0 TO 7);
END COMPONENT;

COMPONENT DECO_7_SEG IS
PORT ( IND_DEC: IN INTEGER RANGE 0 TO 7;
DISPLAY_7_SEG: OUT BIT_VECTOR (6 DOWNTO 0));
END COMPONENT;

BEGIN

CHIP1: DIV_CLK PORT MAP(IN_CLK=> CLK, OUT_CLK=>AUX_CLK_TO_FSM);
CHIP2: FMS_ESTPROJ PORT MAP (IN_CLK=> AUX_CLK_TO_FSM, C1=>SAI_C1, C2=>SAI_C2, C3=>SAI_C3, S1=>ENT_S1, S2=>ENT_S2);
CHIP3: DECO_7_SEG PORT MAP(IND_DEC=>AUX_FMS_TO_DEC, DISPLAY_7_SEG=>DISPLAY_0);
END ONE;


ENTITY FMS_ESTPROJ IS 
PORT(IN_CLK,S1,S2: IN BIT;
C1, C2, C3: OUT BIT;
DISPLAY_7_SEG: OUT INTEGER RANGE 0 TO 7);
END FMS_ESTPROJ;

ARCHITECTURE ONE OF FMS_ESTPROJ IS
TYPE STATE IS (ESTADO_H1,ESTADO_GB,ESTADO_H2,ESTADO_PA,ESTADO_H3,ESTADO_H4,ESTADO_H5,ESTADO_GP);
SIGNAL AUX: STATE;
BEGIN
PROCESS(IN_CLK)
BEGIN
IF (IN_CLK'EVENT)AND(IN_CLK='1') THEN
	CASE AUX IS
	WHEN ESTADO_GP =>
	IF (S1='0' AND S2='1') THEN
	AUX <= ESTADO_H1;
	ELSIF (S1='0' AND S2='0') THEN
	AUX <= ESTADO_H4;
	ELSE 
	AUX <= ESTADO_GP;
	END IF;
	
	WHEN ESTADO_H1 => 
	AUX <= ESTADO_GB;

	WHEN ESTADO_H4 =>
	AUX <= ESTADO_PA;

	WHEN ESTADO_GB =>
	IF (S1='0' AND S2='0') THEN
	AUX <= ESTADO_H2;
	ELSIF (S1='1') THEN
	AUX <= ESTADO_H5;
	ELSE 
	AUX <= ESTADO_GB;
	END IF;
	
	WHEN ESTADO_H2 =>
	AUX<= ESTADO_PA;
	
	WHEN ESTADO_PA =>
	IF (S1='1') THEN
	AUX<= ESTADO_H3;
	ELSE 
	AUX <= ESTADO_PA;
	END IF;
	
	WHEN ESTADO_H3 =>
	AUX <= ESTADO_GP;
	
	WHEN ESTADO_H5 =>
	AUX <= ESTADO_GP;
	
END CASE;
END IF;
END PROCESS;
	
WITH AUX SELECT
	C1<= '1' WHEN ESTADO_GP,
		  '1' WHEN ESTADO_H1,
		  '1' WHEN ESTADO_H4,
		  '0' WHEN OTHERS;
		  
WITH AUX SELECT
   C2<= '1' WHEN ESTADO_H5,
		  '1' WHEN ESTADO_H2,
		  '1' WHEN ESTADO_GB,
		  '0' WHEN OTHERS;
		  
WITH AUX SELECT  
   C3<= '1' WHEN ESTADO_H1,
		  '1' WHEN ESTADO_H4,
		  '1' WHEN ESTADO_GP,
		  '0' WHEN OTHERS;	
		
WITH AUX SELECT
DISPLAY_7_SEG<=   2 	WHEN ESTADO_GB,
						0	WHEN ESTADO_GP, 
						5	WHEN ESTADO_PA,	 
						1	WHEN ESTADO_H1,
						4	WHEN ESTADO_H2,	 
						6	WHEN ESTADO_H3,
						7	WHEN ESTADO_H4, 
						3	WHEN ESTADO_H5;		

END ONE;

		  
ENTITY DIV_CLK IS
PORT(IN_CLK: IN BIT;
OUT_CLK: OUT BIT);
END DIV_CLK;

ARCHITECTURE ONE OF DIV_CLK IS
SIGNAL X: BIT;
SIGNAL Y: INTEGER RANGE 0 TO 4999999:=0;
BEGIN
PROCESS(IN_CLK)
BEGIN
IF (IN_CLK 'EVENT) AND (IN_CLK='1') THEN
	IF Y= 4999999 THEN
	Y<=0;
	X<=NOT (X);
	ELSE
	Y<=Y+1;
	END IF;
END IF;
END PROCESS;
OUT_CLK<=X;
END ONE;

ENTITY DECO_7_SEG IS
PORT ( IND_DEC: IN INTEGER RANGE 0 TO 7;
DISPLAY_7_SEG: OUT BIT_VECTOR (6 DOWNTO 0));
END DECO_7_SEG; 

ARCHITECTURE ONE OF DECO_7_SEG IS
BEGIN
WITH IND_DEC SELECT 
	DISPLAY_7_SEG <=  "0011000" WHEN 0,
							"1001111" WHEN 1,
							"1100000" WHEN 2,
							"0100100" WHEN 3,
							"0010010" WHEN 4,
							"0001000" WHEN 5,
							"0000110" WHEN 6,
							"1001100" WHEN 7;
							
END ONE;			  