ENTITY PRINCIPAL IS
PORT(CLK: IN BIT;
DISPLAY_O: OUT BIT_VECTOR (6 DOWNTO 0);
DISPLAY_1: OUT BIT_VECTOR (6 DOWNTO 0);
DISPLAY_2: OUT BIT_VECTOR (6 DOWNTO 0);
DISPLAY_3: OUT BIT_VECTOR (6 DOWNTO 0);
DISPLAY_4: OUT BIT_VECTOR (6 DOWNTO 0);
DISPLAY_5: OUT BIT_VECTOR (6 DOWNTO 0);
--DISPLAY_6: OUT BIT_VECTOR (6 DOWNTO 0);

TESTE: OUT BIT);
END PRINCIPAL;

ARCHITECTURE ONE OF PRINCIPAL IS  --DECLARA VARIASVEIS DAS INTELIGACOES
SIGNAL AUX: BIT;
SIGNAL DSEG:BIT; -- DESENA DE SEGUNDO
SIGNAL UMIN:BIT; -- UNIDADE DE MINUTO
SIGNAL DMIN:BIT; -- DESENA DE MINUTO	
SIGNAL UHOR:BIT; -- UNIDADE DE HORA
SIGNAL DHOR:BIT; -- DESENA DE HORA
SIGNAL VAICOMDEUS:BIT; -- DECIDIR O USO
SIGNAL AUX_1: INTEGER RANGE 0 TO 9;
SIGNAL AUX_DSEC: INTEGER RANGE 0 TO 5;
SIGNAL AUX_UMIN: INTEGER RANGE 0 TO 9;
SIGNAL AUX_DMIN: INTEGER RANGE 0 TO 9;
SIGNAL AUX_UHOR: INTEGER RANGE 0 TO 9;
SIGNAL AUX_DHOR: INTEGER RANGE 0 TO 9;


COMPONENT DIV_CLK IS
PORT(IN_CLK:IN BIT;
OUT_CLK: OUT BIT);
END COMPONENT;

COMPONENT CONT_9 IS
PORT(IN_CLK, RESET: IN BIT;
SAIDA: OUT INTEGER RANGE 0 TO 9;
COUT:OUT BIT);
END COMPONENT;

COMPONENT DECODIFICADOR_7SEG IS
PORT( DISPLAY: OUT BIT_VECTOR(6 DOWNTO 0);
IN_DEC: IN INTEGER RANGE 0 TO 9);
END COMPONENT;

COMPONENT CONT_5 IS
PORT(IN_CLK, RESET: IN BIT;
SAIDA: OUT INTEGER RANGE 0 TO 5;
COUT:OUT BIT);
END COMPONENT;


BEGIN
CHIP1: DIV_CLK PORT MAP(IN_CLK=> CLK, OUT_CLK=> AUX); -- DIVISO DE CLOCK
CHIP2: CONT_9 PORT MAP (IN_CLK=> AUX, RESET=>'0',SAIDA=>AUX_1,COUT=>DSEG); -- CONTADOR DO USEC
CHIP3: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_O,IN_DEC=> AUX_1); -- DISPLAY DA UNIDADE USEC
CHIP4: CONT_5 PORT MAP(IN_CLK=> DSEG,RESET=>'0', SAIDA=>AUX_DSEC,COUT=>UMIN); -- CONTADOR DO DSEC
CHIP5: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_1,IN_DEC=> AUX_DSEC); -- DISPLAY DSEC
CHIP6: CONT_9 PORT MAP (IN_CLK=> UMIN, RESET=>'0',SAIDA=>AUX_UMIN,COUT=>DMIN); -- CONTADOR DO UMIN
CHIP7: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_2,IN_DEC=> AUX_UMIN); -- DISPLAY UMIN
CHIP8: CONT_5 PORT MAP(IN_CLK=> DMIN,RESET=>'0', SAIDA=>AUX_DMIN,COUT=>UHOR); -- CONTADOR DO DMIN
CHIP9: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_3,IN_DEC=> AUX_DMIN); -- DISPLAY DMIN
CHIP10: CONT_9 PORT MAP (IN_CLK=> UHOR, RESET=>'0',SAIDA=>AUX_UHOR,COUT=>DHOR); -- CONTADOR DO UHOR
CHIP11: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_4,IN_DEC=> AUX_UHOR); -- DISPLAY UHOR
CHIP12: CONT_9 PORT MAP (IN_CLK=> DHOR, RESET=>'0',SAIDA=>AUX_DHOR,COUT=>VAICOMDEUS); -- CONTADOR DO DHOR
CHIP13: DECODIFICADOR_7SEG PORT MAP(DISPLAY=>DISPLAY_5,IN_DEC=> AUX_DHOR); -- DISPLAY DHOR

END ONE;

ENTITY DIV_CLK IS
PORT (in_clk: IN bit;
out_clk: OUT bit);
END DIV_CLK;

ARCHITECTURE master OF DIV_CLK IS
SIGNAL X:bit;
SIGNAL y: integer range 0 to 3999:=0;
--SIGNAL y: integer range 0 to 4999999:=0; ORIGINAL
BEGIN
PROCESS (in_clk)
BEGIN
if (in_clk 'event) and (in_clk='1') then

--if y=4999999 then ORIGINAL
If y=3999 then 
	y<=0;
	x<= not x;
	else
	y<=y+1;
end if;
end if;
end process;
out_clk<=x;
END master;

ENTITY CONT_9 IS
PORT (IN_CLK, RESET: IN BIT;
SAIDA: OUT INTEGER RANGE 0 TO 9;
COUT: OUT BIT);
END CONT_9;

-- CONTADOR DE UNODADE DE SEGUNDO E MINUTO E HORA

ARCHITECTURE MASTER OF CONT_9 IS
SIGNAL AUX_1: BIT;
SIGNAL AUX_2: INTEGER RANGE 0 TO 9;
BEGIN
PROCESS(IN_CLK)
BEGIN
IF RESET='1' THEN
AUX_2<=0;
AUX_1<='0';
ELSIF (IN_CLK'EVENT)AND(IN_CLK='1')THEN
	IF AUX_2=9 THEN
	AUX_2<=0;
   AUX_1<='1';
	ELSE
	AUX_1<='0';
	AUX_2<=AUX_2+1;
	END IF;
END IF;
END PROCESS;
SAIDA<= AUX_2;
COUT<=AUX_1;
END MASTER;

-- DECODIFICADOR DO DISPLAY

ENTITY DECODIFICADOR_7SEG IS
PORT ( DISPLAY: OUT BIT_VECTOR(6 DOWNTO 0);
IN_DEC: IN INTEGER RANGE 0 TO 9);
END DECODIFICADOR_7SEG;

ARCHITECTURE ONE OF DECODIFICADOR_7SEG IS
BEGIN
WITH IN_DEC SELECT
    DISPLAY<=  "0000001" WHEN 0,
					"1001111" WHEN 1,
					"0010010" WHEN 2,
					"0000110" WHEN 3,
					"1001100" WHEN 4,
					"0100100" WHEN 5,
					"0100000" WHEN 6,
					"0001111" WHEN 7,
					"0000000" WHEN 8,
					"0000100" WHEN 9,
					"1111111" WHEN OTHERS;
	 
			  
END ONE;

-- CONTADOR DAS DEZENAS DE SEGUNDOS E MINUTOS

ENTITY CONT_5 IS
PORT (IN_CLK, RESET: IN BIT;
SAIDA: OUT INTEGER RANGE 0 TO 5;
COUT: OUT BIT);
END CONT_5;

ARCHITECTURE MASTER OF CONT_5 IS
SIGNAL AUX_1: BIT;
SIGNAL AUX_2: INTEGER RANGE 0 TO 5;
BEGIN
PROCESS(IN_CLK)
BEGIN
IF RESET='1' THEN
AUX_2<=0;
AUX_1<='0';
ELSIF (IN_CLK'EVENT)AND(IN_CLK='1')THEN
	IF AUX_2=5 THEN
	AUX_2<=0;
   AUX_1<='1';
	ELSE
	AUX_1<='0';
	AUX_2<=AUX_2+1;
	END IF;
END IF;
END PROCESS;
SAIDA<= AUX_2;
COUT<=AUX_1;
END MASTER;


