ENTITY SUBTRATOR IS
PORT(A,B, TE: IN BIT;
S, TS: OUT BIT);
END SUBTRATOR;

ARCHITECTURE ONE OF SUBTRATOR IS 
SIGNAL X: BIT_VECTOR(2 DOWNTO 0);
BEGIN 
X<= A&B&TE;
WITH X SELECT 
   S<= '0' WHEN "000",
	    '1' WHEN "001",
		 '1' WHEN "010",
		 '0' WHEN "011",
		 '1' WHEN "100",
		 '0' WHEN "101",
		 '0' WHEN "110",
		 '1' WHEN "111";
WITH X SELECT 
  TS<= '0' WHEN "000",
	    '1' WHEN "001",
		 '1' WHEN "010",
		 '1' WHEN "011",
		 '0' WHEN "100",
		 '0' WHEN "101",
		 '0' WHEN "110",
		 '1' WHEN "111";
END ONE;

